hello raghavenndra